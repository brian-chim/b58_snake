module game(SW, KEY, CLOCK_50, HEX7, HEX6, HEX5, HEX4, HEX3, HEX2, HEX1, HEX0)
  input KEY[3:2];
  input CLOCK_50;
  input SW[17:0];
  output [6:0] HEX7, HEX6, HEX5, HEX4, HEX3, HEX2, HEX1, HEX0;
  
endmodule


module snake()

endmodule

module tron()

endmodule
