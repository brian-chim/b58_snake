module game(SW, KEY
  input KEY[3:2]

endmodule


module snake

endmodule

module tron

endmodule
